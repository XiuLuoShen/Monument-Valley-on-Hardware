module vga_test(
	input [3:0] KEY,
	input [9:0] SW,
	input CLOCK_50,
	output	[9:0] VGA_R, VGA_G, VGA_B,
	output 	VGA_HS, VGA_VS, VGA_BLANK, VGA_SYNC, VGA_CLK
	);
	
	wire resetn = KEY[0];
	wire ld_dir = ~KEY[1];
	wire move = ~KEY[2];
	wire resetnMonitor = KEY[3];
	wire clear = SW[3];
	wire plot;
	wire [8:0] X;
	wire [7:0] Y;
	wire [2:0] color;
	wire [1:0] dir = SW[1:0];
	
	spriteFSM sprite(
		.clock(CLOCK_50),
		.resetn(resetn),
		.move(move),
		.ld_dir(ld_dir),
		.dir(dir),
		.clear(clear),
		.plot(plot),
		.color(color),
		.xCoord(X),
		.yCoord(Y)
		);
	
	
	vga_adapter display(
		.resetn(resetnMonitor),
		.clock(CLOCK_50),
		.colour(color),
		.x(X),
		.y(Y),
		.plot(plot),
		/* Signals for the DAC to drive the monitor. */
		.VGA_R(VGA_R),
		.VGA_G(VGA_G),
		.VGA_B(VGA_B),
		.VGA_HS(VGA_HS),
		.VGA_VS(VGA_VS),
		.VGA_BLANK(VGA_BLANK),
		.VGA_SYNC(VGA_SYNC),
		.VGA_CLK(VGA_CLK)
	);
	
	defparam display.RESOLUTION = "320x240";
	defparam display.MONOCHROME = "FALSE";
	defparam display.BITS_PER_COLOUR_CHANNEL = 1;
	defparam display.BACKGROUND_IMAGE = "image.colour.mif";
	defparam display.USING_DE1 = "TRUE";
	
endmodule